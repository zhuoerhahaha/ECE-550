module negateb(bin, bout);
	input[31:0] bin;
	output[31:0] bout;
	
	not(bout[0], bin[0]);
	not(bout[1], bin[1]);
	not(bout[2], bin[2]);
	not(bout[3], bin[3]);
	not(bout[4], bin[4]);
	not(bout[5], bin[5]);
	not(bout[6], bin[6]);
	not(bout[7], bin[7]);
	not(bout[8], bin[8]);
	not(bout[9], bin[9]);
	not(bout[10], bin[10]);
	not(bout[11], bin[11]);
	not(bout[12], bin[12]);
	not(bout[13], bin[13]);
	not(bout[14], bin[14]);
	not(bout[15], bin[15]);
	not(bout[16], bin[16]);
	not(bout[17], bin[17]);
	not(bout[18], bin[18]);
	not(bout[19], bin[19]);
	not(bout[20], bin[20]);
	not(bout[21], bin[21]);
	not(bout[22], bin[22]);
	not(bout[23], bin[23]);
	not(bout[24], bin[24]);
	not(bout[25], bin[25]);
	not(bout[26], bin[26]);
	not(bout[27], bin[27]);
	not(bout[28], bin[28]);
	not(bout[29], bin[29]);
	not(bout[30], bin[30]);
	not(bout[31], bin[31]);

	
endmodule
	