module bit_And(ina, inb, out);
	input[31:0] ina, inb;
	output[31:0] out;
	and(out[0], ina[0], inb[0]);
	and(out[1], ina[1], inb[1]);
	and(out[2], ina[2], inb[2]);
	and(out[3], ina[3], inb[3]);
	and(out[4], ina[4], inb[4]);
	and(out[5], ina[5], inb[5]);
	and(out[6], ina[6], inb[6]);
	and(out[7], ina[7], inb[7]);
	and(out[8], ina[8], inb[8]);
	and(out[9], ina[9], inb[9]);
	and(out[10], ina[10], inb[10]);
	and(out[11], ina[11], inb[11]);
	and(out[12], ina[12], inb[12]);
	and(out[13], ina[13], inb[13]);
	and(out[14], ina[14], inb[14]);
	and(out[15], ina[15], inb[15]);
	and(out[16], ina[16], inb[16]);
	and(out[17], ina[17], inb[17]);
	and(out[18], ina[18], inb[18]);
	and(out[19], ina[19], inb[19]);
	and(out[20], ina[20], inb[20]);
	and(out[21], ina[21], inb[21]);
	and(out[22], ina[22], inb[22]);
	and(out[23], ina[23], inb[23]);
	and(out[24], ina[24], inb[24]);
	and(out[25], ina[25], inb[25]);
	and(out[26], ina[26], inb[26]);
	and(out[27], ina[27], inb[27]);
	and(out[28], ina[28], inb[28]);
	and(out[29], ina[29], inb[29]);
	and(out[30], ina[30], inb[30]);
	and(out[31], ina[31], inb[31]);
endmodule
	
	