module multipleAND(in, out, en);
	input[31:0] in;
	input en;
	output[31:0] out;
	
	
	and and0(out[0], in[0], en);
	and and1(out[1], in[1], en);
	and and2(out[2], in[2], en);
	and and3(out[3], in[3], en);
	and and4(out[4], in[4], en);
	and and5(out[5], in[5], en);
	and and6(out[6], in[6], en);
	and and7(out[7], in[7], en);
	and and8(out[8], in[8], en);
	and and9(out[9], in[9], en);
	and and10(out[10], in[10], en);
	and and11(out[11], in[11], en);
	and and12(out[12], in[12], en);
	and and13(out[13], in[13], en);
	and and14(out[14], in[14], en);
	and and15(out[15], in[15], en);
	and and16(out[16], in[16], en);
	and and17(out[17], in[17], en);
	and and18(out[18], in[18], en);
	and and19(out[19], in[19], en);
	and and20(out[20], in[20], en);
	and and21(out[21], in[21], en);
	and and22(out[22], in[22], en);
	and and23(out[23], in[23], en);
	and and24(out[24], in[24], en);
	and and25(out[25], in[25], en);
	and and26(out[26], in[26], en);
	and and27(out[27], in[27], en);
	and and28(out[28], in[28], en);
	and and29(out[29], in[29], en);
	and and30(out[30], in[30], en);
	and and31(out[31], in[31], en);
endmodule