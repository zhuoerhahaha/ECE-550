module bit_Or(ina, inb, out);
	input[31:0] ina, inb;
	output[31:0] out;
	or(out[0], ina[0], inb[0]);
	or(out[1], ina[1], inb[1]);
	or(out[2], ina[2], inb[2]);
	or(out[3], ina[3], inb[3]);
	or(out[4], ina[4], inb[4]);
	or(out[5], ina[5], inb[5]);
	or(out[6], ina[6], inb[6]);
	or(out[7], ina[7], inb[7]);
	or(out[8], ina[8], inb[8]);
	or(out[9], ina[9], inb[9]);
	or(out[10], ina[10], inb[10]);
	or(out[11], ina[11], inb[11]);
	or(out[12], ina[12], inb[12]);
	or(out[13], ina[13], inb[13]);
	or(out[14], ina[14], inb[14]);
	or(out[15], ina[15], inb[15]);
	or(out[16], ina[16], inb[16]);
	or(out[17], ina[17], inb[17]);
	or(out[18], ina[18], inb[18]);
	or(out[19], ina[19], inb[19]);
	or(out[20], ina[20], inb[20]);
	or(out[21], ina[21], inb[21]);
	or(out[22], ina[22], inb[22]);
	or(out[23], ina[23], inb[23]);
	or(out[24], ina[24], inb[24]);
	or(out[25], ina[25], inb[25]);
	or(out[26], ina[26], inb[26]);
	or(out[27], ina[27], inb[27]);
	or(out[28], ina[28], inb[28]);
	or(out[29], ina[29], inb[29]);
	or(out[30], ina[30], inb[30]);
	or(out[31], ina[31], inb[31]);
endmodule