module right_shift(in, shiftamout, out);
	input[31:0] in;
	input[4:0] shiftamout;
	
	output[31:0] out;
	
endmodule
